module HISTOGRAM_1CELL (

	input iClk,
	input [7:0] iPX11, iPX12, iPX13, iPX14, iPX15, iPX16, iPX17, iPX18, iPX19, iPX1_10, 
	input [7:0] iPX21, iPX22, iPX23, iPX24, iPX25, iPX26, iPX27, iPX28, iPX29, iPX2_10, 
	input [7:0] iPX31, iPX32, iPX33, iPX34, iPX35, iPX36, iPX37, iPX38, iPX39, iPX3_10, 
	input [7:0] iPX41, iPX42, iPX43, iPX44, iPX45, iPX46, iPX47, iPX48, iPX49, iPX4_10, 
	input [7:0] iPX51, iPX52, iPX53, iPX54, iPX55, iPX56, iPX57, iPX58, iPX59, iPX5_10, 
	input [7:0] iPX61, iPX62, iPX63, iPX64, iPX65, iPX66, iPX67, iPX68, iPX69, iPX6_10, 
	input [7:0] iPX71, iPX72, iPX73, iPX74, iPX75, iPX76, iPX77, iPX78, iPX79, iPX7_10, 
	input [7:0] iPX81, iPX82, iPX83, iPX84, iPX85, iPX86, iPX87, iPX88, iPX89, iPX8_10, 
	input [7:0] iPX91, iPX92, iPX93, iPX94, iPX95, iPX96, iPX97, iPX98, iPX99, iPX9_10, 
	input [7:0] iPX10_1, iPX10_2, iPX10_3, iPX10_4, iPX10_5, iPX10_6, iPX10_7, iPX10_8, iPX10_9, iPX10_10,
	
	output [31:0] oBIN1, oBIN2, oBIN3, oBIN4, oBIN5, oBIN6, oBIN7, oBIN8, oBIN9
);


	// 64 32-bits output magnitude values.
	wire [31:0] oMAG11, oMAG12, oMAG13, oMAG14, oMAG15, oMAG16, oMAG17, oMAG18; 
	wire [31:0] oMAG21, oMAG22, oMAG23, oMAG24, oMAG25, oMAG26, oMAG27, oMAG28; 
	wire [31:0] oMAG31, oMAG32, oMAG33, oMAG34, oMAG35, oMAG36, oMAG37, oMAG38; 
	wire [31:0] oMAG41, oMAG42, oMAG43, oMAG44, oMAG45, oMAG46, oMAG47, oMAG48; 
	wire [31:0] oMAG51, oMAG52, oMAG53, oMAG54, oMAG55, oMAG56, oMAG57, oMAG58; 
	wire [31:0] oMAG61, oMAG62, oMAG63, oMAG64, oMAG65, oMAG66, oMAG67, oMAG68; 
	wire [31:0] oMAG71, oMAG72, oMAG73, oMAG74, oMAG75, oMAG76, oMAG77, oMAG78; 
	wire [31:0] oMAG81, oMAG82, oMAG83, oMAG84, oMAG85, oMAG86, oMAG87, oMAG88;  

	// 64 32-bits output angle values.
	wire [31:0] oAGL11, oAGL12, oAGL13, oAGL14, oAGL15, oAGL16, oAGL17, oAGL18; 
	wire [31:0] oAGL21, oAGL22, oAGL23, oAGL24, oAGL25, oAGL26, oAGL27, oAGL28; 
	wire [31:0] oAGL31, oAGL32, oAGL33, oAGL34, oAGL35, oAGL36, oAGL37, oAGL38; 
	wire [31:0] oAGL41, oAGL42, oAGL43, oAGL44, oAGL45, oAGL46, oAGL47, oAGL48; 
	wire [31:0] oAGL51, oAGL52, oAGL53, oAGL54, oAGL55, oAGL56, oAGL57, oAGL58; 
	wire [31:0] oAGL61, oAGL62, oAGL63, oAGL64, oAGL65, oAGL66, oAGL67, oAGL68; 
	wire [31:0] oAGL71, oAGL72, oAGL73, oAGL74, oAGL75, oAGL76, oAGL77, oAGL78; 
	wire [31:0] oAGL81, oAGL82, oAGL83, oAGL84, oAGL85, oAGL86, oAGL87, oAGL88;
	
	
	
	GRADIENT_1CELL GRADIENT_1CELL(
	
		.iClk(iClk),
		// We need 10x10 input pixels for computing gradient of 64 pixels (including 36 pixels on the border).
		// Input values are 8-bits values. 
		.iPX11(iPX11), .iPX12(iPX12), .iPX13(iPX13), .iPX14(iPX14), .iPX15(iPX15), .iPX16(iPX16), .iPX17(iPX17), .iPX18(iPX18), .iPX19(iPX19), .iPX1_10(iPX1_10), 
		.iPX21(iPX21), .iPX22(iPX22), .iPX23(iPX23), .iPX24(iPX24), .iPX25(iPX25), .iPX26(iPX26), .iPX27(iPX27), .iPX28(iPX28), .iPX29(iPX29), .iPX2_10(iPX2_10), 
		.iPX31(iPX31), .iPX32(iPX32), .iPX33(iPX33), .iPX34(iPX34), .iPX35(iPX35), .iPX36(iPX36), .iPX37(iPX37), .iPX38(iPX38), .iPX39(iPX39), .iPX3_10(iPX3_10), 
		.iPX41(iPX41), .iPX42(iPX42), .iPX43(iPX43), .iPX44(iPX44), .iPX45(iPX45), .iPX46(iPX46), .iPX47(iPX47), .iPX48(iPX48), .iPX49(iPX49), .iPX4_10(iPX4_10), 
		.iPX51(iPX51), .iPX52(iPX52), .iPX53(iPX53), .iPX54(iPX54), .iPX55(iPX55), .iPX56(iPX56), .iPX57(iPX57), .iPX58(iPX58), .iPX59(iPX59), .iPX5_10(iPX5_10), 
		.iPX61(iPX61), .iPX62(iPX62), .iPX63(iPX63), .iPX64(iPX64), .iPX65(iPX65), .iPX66(iPX66), .iPX67(iPX67), .iPX68(iPX68), .iPX69(iPX69), .iPX6_10(iPX6_10), 
		.iPX71(iPX71), .iPX72(iPX72), .iPX73(iPX73), .iPX74(iPX74), .iPX75(iPX75), .iPX76(iPX76), .iPX77(iPX77), .iPX78(iPX78), .iPX79(iPX79), .iPX7_10(iPX7_10), 
		.iPX81(iPX81), .iPX82(iPX82), .iPX83(iPX83), .iPX84(iPX84), .iPX85(iPX85), .iPX86(iPX86), .iPX87(iPX87), .iPX88(iPX88), .iPX89(iPX89), .iPX8_10(iPX8_10), 
		.iPX91(iPX91), .iPX92(iPX92), .iPX93(iPX93), .iPX94(iPX94), .iPX95(iPX95), .iPX96(iPX96), .iPX97(iPX97), .iPX98(iPX98), .iPX99(iPX99), .iPX9_10(iPX9_10), 
		.iPX10_1(iPX10_1), .iPX10_2(iPX10_2), .iPX10_3(iPX10_3), .iPX10_4(iPX10_4), .iPX10_5(iPX10_5), .iPX10_6(iPX10_6), .iPX10_7(iPX10_7), .iPX10_8(iPX10_8), .iPX10_9(iPX10_9), .iPX10_10(iPX10_10), 

		// We will have 64 output gradient values
		// Each output gradient value includes a magnitude value and a angle value in floating-point index.
		// Totally, we will have 128 32-bits output values.

		// 64 32-bits output magnitude values.
		.oMAG11(oMAG11), .oMAG12(oMAG12), .oMAG13(oMAG13), .oMAG14(oMAG14), .oMAG15(oMAG15), .oMAG16(oMAG16), .oMAG17(oMAG17), .oMAG18(oMAG18), 
		.oMAG21(oMAG21), .oMAG22(oMAG22), .oMAG23(oMAG23), .oMAG24(oMAG24), .oMAG25(oMAG25), .oMAG26(oMAG26), .oMAG27(oMAG27), .oMAG28(oMAG28), 
		.oMAG31(oMAG31), .oMAG32(oMAG32), .oMAG33(oMAG33), .oMAG34(oMAG34), .oMAG35(oMAG35), .oMAG36(oMAG36), .oMAG37(oMAG37), .oMAG38(oMAG38), 
		.oMAG41(oMAG41), .oMAG42(oMAG42), .oMAG43(oMAG43), .oMAG44(oMAG44), .oMAG45(oMAG45), .oMAG46(oMAG46), .oMAG47(oMAG47), .oMAG48(oMAG48), 
		.oMAG51(oMAG51), .oMAG52(oMAG52), .oMAG53(oMAG53), .oMAG54(oMAG54), .oMAG55(oMAG55), .oMAG56(oMAG56), .oMAG57(oMAG57), .oMAG58(oMAG58), 
		.oMAG61(oMAG61), .oMAG62(oMAG62), .oMAG63(oMAG63), .oMAG64(oMAG64), .oMAG65(oMAG65), .oMAG66(oMAG66), .oMAG67(oMAG67), .oMAG68(oMAG68), 
		.oMAG71(oMAG71), .oMAG72(oMAG72), .oMAG73(oMAG73), .oMAG74(oMAG74), .oMAG75(oMAG75), .oMAG76(oMAG76), .oMAG77(oMAG77), .oMAG78(oMAG78), 
		.oMAG81(oMAG81), .oMAG82(oMAG82), .oMAG83(oMAG83), .oMAG84(oMAG84), .oMAG85(oMAG85), .oMAG86(oMAG86), .oMAG87(oMAG87), .oMAG88(oMAG88),  

		// 64 32-bits output angle values.
		.oAGL11(oAGL11), .oAGL12(oAGL12), .oAGL13(oAGL13), .oAGL14(oAGL14), .oAGL15(oAGL15), .oAGL16(oAGL16), .oAGL17(oAGL17), .oAGL18(oAGL18), 
		.oAGL21(oAGL21), .oAGL22(oAGL22), .oAGL23(oAGL23), .oAGL24(oAGL24), .oAGL25(oAGL25), .oAGL26(oAGL26), .oAGL27(oAGL27), .oAGL28(oAGL28), 
		.oAGL31(oAGL31), .oAGL32(oAGL32), .oAGL33(oAGL33), .oAGL34(oAGL34), .oAGL35(oAGL35), .oAGL36(oAGL36), .oAGL37(oAGL37), .oAGL38(oAGL38), 
		.oAGL41(oAGL41), .oAGL42(oAGL42), .oAGL43(oAGL43), .oAGL44(oAGL44), .oAGL45(oAGL45), .oAGL46(oAGL46), .oAGL47(oAGL47), .oAGL48(oAGL48), 
		.oAGL51(oAGL51), .oAGL52(oAGL52), .oAGL53(oAGL53), .oAGL54(oAGL54), .oAGL55(oAGL55), .oAGL56(oAGL56), .oAGL57(oAGL57), .oAGL58(oAGL58), 
		.oAGL61(oAGL61), .oAGL62(oAGL62), .oAGL63(oAGL63), .oAGL64(oAGL64), .oAGL65(oAGL65), .oAGL66(oAGL66), .oAGL67(oAGL67), .oAGL68(oAGL68), 
		.oAGL71(oAGL71), .oAGL72(oAGL72), .oAGL73(oAGL73), .oAGL74(oAGL74), .oAGL75(oAGL75), .oAGL76(oAGL76), .oAGL77(oAGL77), .oAGL78(oAGL78), 
		.oAGL81(oAGL81), .oAGL82(oAGL82), .oAGL83(oAGL83), .oAGL84(oAGL84), .oAGL85(oAGL85), .oAGL86(oAGL86), .oAGL87(oAGL87), .oAGL88(oAGL88)

		);
		
	GETHISTOGRAM_1CELL GETHISTOGRAM_1CELL(

  .iClk(iClk),
  .iMAG11(oMAG11), .iMAG12(oMAG12), .iMAG13(oMAG13), .iMAG14(oMAG14), .iMAG15(oMAG15), .iMAG16(oMAG16), .iMAG17(oMAG17), .iMAG18(oMAG18), 
  .iMAG21(oMAG21), .iMAG22(oMAG22), .iMAG23(oMAG23), .iMAG24(oMAG24), .iMAG25(oMAG25), .iMAG26(oMAG26), .iMAG27(oMAG27), .iMAG28(oMAG28), 
  .iMAG31(oMAG31), .iMAG32(oMAG32), .iMAG33(oMAG33), .iMAG34(oMAG34), .iMAG35(oMAG35), .iMAG36(oMAG36), .iMAG37(oMAG37), .iMAG38(oMAG38), 
  .iMAG41(oMAG41), .iMAG42(oMAG42), .iMAG43(oMAG43), .iMAG44(oMAG44), .iMAG45(oMAG45), .iMAG46(oMAG46), .iMAG47(oMAG47), .iMAG48(oMAG48), 
  .iMAG51(oMAG51), .iMAG52(oMAG52), .iMAG53(oMAG53), .iMAG54(oMAG54), .iMAG55(oMAG55), .iMAG56(oMAG56), .iMAG57(oMAG57), .iMAG58(oMAG58), 
  .iMAG61(oMAG61), .iMAG62(oMAG62), .iMAG63(oMAG63), .iMAG64(oMAG64), .iMAG65(oMAG64), .iMAG66(oMAG66), .iMAG67(oMAG67), .iMAG68(oMAG68), 
  .iMAG71(oMAG71), .iMAG72(oMAG72), .iMAG73(oMAG73), .iMAG74(oMAG74), .iMAG75(oMAG75), .iMAG76(oMAG76), .iMAG77(oMAG77), .iMAG78(oMAG78), 
  .iMAG81(oMAG81), .iMAG82(oMAG82), .iMAG83(oMAG83), .iMAG84(oMAG84), .iMAG85(oMAG85), .iMAG86(oMAG86), .iMAG87(oMAG87), .iMAG88(oMAG88), 
  
  .iAGL11(oAGL11), .iAGL12(oAGL12), .iAGL13(oAGL13), .iAGL14(oAGL14), .iAGL15(oAGL15), .iAGL16(oAGL16), .iAGL17(oAGL17), .iAGL18(oAGL18), 
  .iAGL21(oAGL21), .iAGL22(oAGL22), .iAGL23(oAGL23), .iAGL24(oAGL24), .iAGL25(oAGL25), .iAGL26(oAGL26), .iAGL27(oAGL27), .iAGL28(oAGL28), 
  .iAGL31(oAGL31), .iAGL32(oAGL32), .iAGL33(oAGL33), .iAGL34(oAGL34), .iAGL35(oAGL35), .iAGL36(oAGL36), .iAGL37(oAGL37), .iAGL38(oAGL38), 
  .iAGL41(oAGL41), .iAGL42(oAGL42), .iAGL43(oAGL43), .iAGL44(oAGL44), .iAGL45(oAGL45), .iAGL46(oAGL46), .iAGL47(oAGL47), .iAGL48(oAGL48), 
  .iAGL51(oAGL51), .iAGL52(oAGL52), .iAGL53(oAGL53), .iAGL54(oAGL54), .iAGL55(oAGL55), .iAGL56(oAGL56), .iAGL57(oAGL57), .iAGL58(oAGL58), 
  .iAGL61(oAGL61), .iAGL62(oAGL62), .iAGL63(oAGL63), .iAGL64(oAGL64), .iAGL65(oAGL65), .iAGL66(oAGL66), .iAGL67(oAGL67), .iAGL68(oAGL68), 
  .iAGL71(oAGL71), .iAGL72(oAGL72), .iAGL73(oAGL73), .iAGL74(oAGL74), .iAGL75(oAGL75), .iAGL76(oAGL76), .iAGL77(oAGL77), .iAGL78(oAGL78), 
  .iAGL81(oAGL81), .iAGL82(oAGL82), .iAGL83(oAGL83), .iAGL84(oAGL84), .iAGL85(oAGL85), .iAGL86(oAGL86), .iAGL87(oAGL87), .iAGL88(oAGL88), 
  
  .oBIN1(oBIN1), .oBIN2(oBIN2), .oBIN3(oBIN3), .oBIN4(oBIN4), .oBIN5(oBIN5), .oBIN6(oBIN6), .oBIN7(oBIN7), .oBIN8(oBIN8), .oBIN9(oBIN9)
  
);

endmodule

